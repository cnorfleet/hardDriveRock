module testbench();
	
endmodule
